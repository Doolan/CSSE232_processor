// Verilog test fixture created from schematic /home/xniccum/projects/csse232/1415a-csse232-niccumas/CSSE232_processor/Components/Processor.sch - Wed Nov  5 16:17:36 2014

`timescale 1ns / 1ps

module Processor_Processor_sch_tb();

// Inputs

// Output

// Bidirs

// Instantiate the UUT
   Processor UUT (
		
   );
// Initialize Inputs
   `ifdef auto_init
       initial begin
   `endif
endmodule
